// acoustic data collection with FPGA

//
// clock counter, enable is active low, after 14 clock cycles, toggle enable
module Datapath(input ); 

endmodule


 