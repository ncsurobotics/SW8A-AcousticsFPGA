// March 11 pool test controller
// submodules: SIPO_Controller, counter, Test_State_Machine

module Test_Controller (
                            input clk,
                            input reset_b
);


endmodule