module top(
    



);

endmodule