module data_buffer();

endmodule