module cross correlator();


endmodule