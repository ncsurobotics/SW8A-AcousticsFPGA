
module header(output wire [800:0] workspace_path);
    assign workspace_path = "C:Users/ilena/Documents/apr-private/fpga/SW8A-AcousticsFPGA";
endmodule