module FFT();

endmodule