

module UART_tb;

endmodule