module UART_tx_datapath #(
    parameter BAUD = 11'868
) (
    
);
    
endmodule