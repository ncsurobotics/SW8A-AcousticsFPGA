module UART();


endmodule